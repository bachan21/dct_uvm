`include "dct_intf.sv"
`include "dct_sequence_item.sv"
`include "sequence_files.sv"
`include "dct_sequence.sv"
`include "dct_sequencer.sv"
`include "dct_driver.sv"
`include "dct_monitor.sv"
`include "dct_agent.sv"
`include "dct_ref_model.sv"
`include "dct_scoreboard.sv"
`include "dct_env.sv"
`include "dct_test.sv"
